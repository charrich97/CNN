module MyDesign
(
//////////////////////////////////////////////////////////////////////////////////
//Clock and Reset Schema
//////////////////////////////////////////////////////////////////////////////////
input               clk                   ,
input               reset_b               ,  

//////////////////////////////////////////////////////////////////////////////////
//Control signals
//////////////////////////////////////////////////////////////////////////////////
input               dut_run               , 
output wire         dut_busy              ,

//////////////////////////////////////////////////////////////////////////////////
//Input and Weight Matrix Addressing
//////////////////////////////////////////////////////////////////////////////////
output wire [11:0]  dut_sram_read_address ,
output wire [11:0]  dut_wmem_read_address ,

//////////////////////////////////////////////////////////////////////////////////
//Input and Weight Matrix Data
//////////////////////////////////////////////////////////////////////////////////
input       [15:0]  sram_dut_read_data    ,
input       [15:0]  wmem_dut_read_data    ,

//////////////////////////////////////////////////////////////////////////////////
//Write Output Signals
//////////////////////////////////////////////////////////////////////////////////
output wire         dut_sram_write_enable , 
output wire [11:0]  dut_sram_write_address,
output wire [15:0]  dut_sram_write_data   
);

//////////////////////////////////////////////////////////////////////////////////
//Interfacing to CNN Device Under Test
//////////////////////////////////////////////////////////////////////////////////
CNN_DUT DUT
(
.go                 (dut_run                ),
.busy               (dut_busy               ),
.clk              	(clk                    ),
.reset              (reset_b                ),
.Write_Address      (dut_sram_write_address ),
.Write_Data         (dut_sram_write_data    ),
.Write_Enable       (dut_sram_write_enable  ),
.Matrix_Address     (dut_sram_read_address  ),
.Read_Matrix_Data   (sram_dut_read_data     ),
.Weight_Address     (dut_wmem_read_address  ),
.Read_Weight_Data   (wmem_dut_read_data     )
);

endmodule
